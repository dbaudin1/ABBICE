* ADA4627 SPICE Macro-model                   
* Description: Amplifier
* Generic Desc: 8/30V, JFET, OP, Low Noise, Low Ib, 1X
* Developed by: HH / ADSJ
* Revision History: 08/10/2012 - Updated to new header style
* 1.0 (07/2009)
* Copyright 2009, 2012 by Analog Devices
*
* Refer to http://www.analog.com/Analog_Root/static/techSupport/designTools/spiceModels/license/spice_general.html for License Statement.  Use of this model
* indicates your acceptance of the terms and provisions in the License Statement.
*
* BEGIN Notes: 
*  CAUTION!!  To aid in convergence, most Spice simulators add a
*  conductance on every node to insure that no node is floating.
*  This is GMIN, and the default value is usually 1E-12. To properly 
*  simulate the low input bias current and low current noise, the 
*  Spice simulator options have to be set to the following:
*  .OPTIONS GMIN=0.01p
*  .OPTIONS ABSTOL=0.01pA
*  .OPTIONS ITL1=500
*  .OPTIONS ITL2=200
*  .OPTIONS ITL4=100
*
* Not Modeled:
*    
* Parameters modeled include: 
*
* END Notes
*
* Node assignments
*                 non-inverting input
*                 |   inverting input
*                 |   |    positive supply
*                 |   |    |    negative supply
*                 |   |    |    |    output
*                 |   |    |    |    |
.SUBCKT ADA4627   1   2   99   50   30
*
* INPUT STAGE
*
Cdiff 1   2  4.7E-12
Cin1  1  50  7.5E-12
Cin2  2  50  7.5E-12
*
R3   5  99    1.478E+03
R4   6  99    1.478E+03
J1   5   2    4   JX
J2   6   7    4   JX
*
I1   4  50    2.70E-03
DI1  4a  4   DX
VI1  4a 50  5.5V
IOS  1   2    0.25E-12
EOS  60  1    POLY(2)  (17,24) (73,98) 110E-6  1  1
EN   7  60    42  0  1
*
EREF 98  0    24  0   1
*
* SECOND STAGE 
*
R5   9  98    4.097E+05
C3   9  98    3.850E-09
G1   98  9    5  6  7.700E-02
V2   99  8    2.86
V3   10 50    2.41;
D1   9   8    DX
D2   10  9    DX
*
* 2nd POLE
*
R13  18 98     1.000E+03
C9   18 98     1.0E-14
G5   98 18     9  24  1E-3
*
* COMMON-MODE GAIN NETWORK 
*
R11  16 17     2.698E-01
R12  17 98     1.326E-04
E3   16 98     POLY(2) 1  98  2  98  0  8.459E-03 8.459E-03
C8   16 17     100E-6
*
* PSRR NETWORK
*
EPSY 98 72 POLY(1) (99,50) 3.350E-03  1.005E-01
CPS3 72 73 1.000E-09
RPS3 72 73 9.947E+05
RPS4 73 98 1.326E+02
*
* VOLTAGE NOISE GENERATOR
*
VN1  41  0    DC 2
DN1  41 42    DEN
DN2  42 43    DEN
VN2  0  43    DC 2
*
* CURRENT NOISE GENERATOR
*
VN3  44  0    DC 2
DN3  44 45    DIN
DN4  45 46    DIN
VN4  0  46    DC 2
*
* CURRENT NOISE GENERATOR
*
VN5  47  0    DC 2
DN5  47 48    DIN
DN6  48 49    DIN
VN6  0  49    DC 2
*
* OUTPUT STAGE
*
R14  24 99     500E3
R15  24 50     500E3
GSY  99 50 POLY(1) (99,50) 4.079E-03 2.985E-06
R16  29 99     100
R17  29 50     100
G6   27 50 18 29  10.0E-3 
G7   28 50 29 18  10.0E-3
G8   29 99  POLY(1)    99 18  1E-16 1.00E-2 
G9   50 29  POLY(1)    18 50  1E-16 1.00E-2
*
V4   25 29     1.99; Isc high side
V5   29 26     2.4
D3   18 25     DX
D4   26 18     DX
*
D5   99 27     DX
D6   99 28     DX
D7   50 27     DY
D8   50 28     DY
F1   29  0     V4  1
F2   0  29     V5  1
L1   29 30a     1E-15
R24  30a 30  1m
*
* MODELS USED
*
.MODEL JX NJF(BETA=3.400E-03  VTO=-1.500  IS=7E-13 RD=1
+ RS=1 CGD=1.5E-12 CGS=1.5E-12 )
*.MODEL JX PJF(BETA=1.4E-3  VTO=-1.000  IS=20E-12 RD=0
*+ RS=0 CGD=3E-12 CGS=3E-12)
.MODEL DX   D(IS=1E-15 RS=0 CJO=1E-12)
.MODEL DY   D(IS=1E-15 BV=50 RS=10 CJO=1E-12)
.MODEL DEN  D(IS=1E-12 RS=1.7E3, KF=6.53E-15 AF=1)
.MODEL DIN  D(IS=1E-12 RS=12090 KF=0 AF=1)
*
.ENDS ADA4627
$




