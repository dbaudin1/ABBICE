* AD8022 Spice Model
* Description: Amplifier
* Generic Desc: Dual high speed low noise amplifier
* Developed by: TRW
* Revision History: 08/10/2012 - Updated to new header style
* 3.0 ( 01/2000)
* Copyright 2000, 2012 by Analog Devices, Inc.
*
* Refer to http://www.analog.com/Analog_Root/static/techSupport/designTools/spiceModels/license/spice_general.html for License Statement.
* Use of this model indicates your acceptance with the terms and provisions in the License Statement
*
* BEGIN Notes:
*
* Not Modeled:
*       distortion is not characterized
*
* Parameters modeled include:
*       open loop gain and phase vs. frequency
*       output clamping voltage and current
*       input common mode range
*       slew rate
*       output currents are reflected to V supplies
*       Vos is static and will not vary
*       step response is modeled at
*
* END Notes
*
* Node assignments
*                   non-inverting input
*                   | inverting input
*                   | | positive supply
*                   | | |  negative supply
*                   | | |  |  output
*                   | | |  |  |
.subckt AD8022      1 2 99 50 23

***** Input stage

Q1 3 4 5 nbjt
Q2 6 1 7 nbjt
Rc1 99 3 118
Rc2 99 6 118
Re1 5 8 31
Re2 8 7 31
I1 8 50 0.6m
D1 9 8 diode
Vdiode 50 9 -.72
Eos 4 2 poly(1) 40 98 2.9m 1

***** Input Error Sources

Cin1 1 98 0.7pF
Cin2 2 98 0.7pF
RinDiff 1 2 20k

****** Gain Stage

Ggain1 10 98 6 3 .00955
Rgain1 10 98 589k
Cgain1 10 98 12pF
Doutclamp1 10 11 diode
Voutclamp1 99 11 2.5
Doutlclamp2 12 10 diode
Voutclamp2 12 50 2.5

****** Reference Stage

Eref1 98 0 poly(2) 99 0 50 0 0 0.5 0.5
Eref2 97 0 poly(2) 1 0 2 0 0 0.5 0.5

***** CMRR Stage

Gcmrr 40 98 98 97 .55e-10
Rc 98 41 1e6
Lc 40 41 8

****** Output Stage

Dout1 10 20 diode
Dout2 21 10 diode
V1 20 22 -0.741
V2 22 21 -0.741
Go1 22 99 99 10 15.823
Go2 50 22 10 50 15.823
Rout1 99 22 .0632
Rout2 22 50 .0632
Vcd 23 22 0

foo1 98 70 vcd 1
Do1 70 71 diode
Do2 72 70 diode
vi1 98 71 0
vi2 72 98 0

Erefq 96 0 23 0 1
Iq 99 50 6.0m
Fq1 99 96 poly(2) vi2 vcd 0 -1 0.5
Fq2 96 50 poly(2) vi1 vcd 0 -1 -0.5


.model diode D(IS=1e-15)
.model nbjt npn(bf=150)
.ends






