* MAX4106 FAMILY MACROMODELS
* -------------------------
* FEATURES:
* 350MHz -3dB Bandwidth
* 15mA Typical Supply Current
* 80mA Output Drive
* 275V/uS Slew Rate
* Available in 8-Pin SO 
*
* PART NUMBER    DESCRIPTION
* ___________    ______________________________
* MAX4106        350MHz, Ultra-Low-Noise Op Amp  
*
*
*   ////////////// MAX4106 MACROMODEL //////////////////
*
*   ====>      REFER TO MAX4106 DATA SHEET       <====
*
* connections:          non-inverting input
*                       |       inverting input
*                       |       |       positive power-supply
*                       |       |       |       negative power-supply
*                       |       |       |       |       output
*                       |       |       |       |       |
* OUTPUT CONNECTS:      1       2       99      50      97
*
* NOTE OFFSET HAS NOT BEEN ADDED TO THIS MODEL 
*
.SUBCKT MAX4106 1 2 99 50 97
****************INPUT STAGE**********************
*
IOS 2 1 50N
I1 4 50 2MA
GIN 2 1 2 1 50E-9
*CIN 1 2 4PF
G16 0 1 106 0 .87E-3
G19 0 2 109 0 .87E-3
****VCCS NOISE INPUT CURRENTS****
G1 5 99 5 99 38.5E-3
G2 6 99 6 99 38.5E-3
vos 1 3 0v
*EOS 1 3 POLY(1) 98 30 0 .63
*               ^       OFFSET VOLTAGE

*****OFFSET VOLTAGE MUST BE 0V TO PERFORM SMALL-SIGNAL ANALYSIS*****
*Vn 3 9 0v
EN 3 9 POLY(1) 103 0 0 .70
Q1 5 2 4 QX
Q2 6 9 4 QX
Dsub 50 99 DX
C4 5 6 6PF
*
*****************NOISE GENERATORS**************
*
***VOLTAGE NOISE GENERATOR***
VN1 101 0 2V
VN2 0 102 2V 
DN1 101 103 D1
DN2 103 102 D1
.MODEL D1 D(KF=10E-15 RS=33)
****CURRENT NOISE GENERATOR + IN****
VN3 104 0 2V
VN4 0 105 2V
DN3 104 106 D2
DN4 106 105 D2
****CURRENT NOISE GENERATOR - IN****
VN5 107 0 2V
VN6 0 108 2V
DN5 107 109 D2
DN6 109 108 D2
.MODEL D2 D(KF=30E-16 RS=20)
*
***************SECOND STAGE******************
IS 99 50 13mA
*         SETS IS ^
****OUTPUT VOLTAGE LIMITING****
V2 99 11 .5
D1 12 11 DX
D2 10 12 DX
V3 10 50 .5
****LEVEL TRANSLATION ****
EH 99 98 99 50 0.5
****GAIN, 1ST POLE****
G3 98 12 5 6 27.1E-3
*27.1
*1ST POLE 21HZ,AVOL 1E6
r4 12 98 6254E3
C3 98 12 2.1E-12
*1.78
*    2.32
**************FREQUENCY SHAPING STAGES********
*
****POLE STAGE****
*G5 98 15 12 98 1E-3 
*G6 98 15 98 15 1E-3
*D13 50 15 DX
*R5 98 15 1E3
*C5 98 15 2.45E-12
*                  ^ POLE AT 65MEGHZ
****COMMON-MODE STAGE****
G11 98 30 4 98 316E-12
G13 30 98 30 98 1E-3
D11 50 30 DX
*
*******************OUTPUT STAGE****************
F6 99 50 VA7 1
F5 99 38 VA8 1
D9 40 38 DX
D10 38 99 DX
VA7 99 40 0
****************
G12 98 32 12 98 1E-3
R15 98 32 1E3
D3 32 36 DX
D4 37 32 DX
V5 35 37 4V
V4 36 35 4V
R16 34 35 30
E1 99 33 99 32 1
VA8 33 34 0V
L 35 96 50P
R17 96 97 20
*
***** MODELS USED ******
.MODEL DX D(IS=1E-15)
.MODEL QX NPN(BF=55.5)
*BF IS SET FOR FOR INPUT BIAS
.ends